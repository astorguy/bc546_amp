.title circuit
.include ./models.sp
.include ./stimulus.sp
.include ./supplies.sp
.include ./load.sp
.include ./dut.sp
.include ./control.sp
.end
